module uart_tfifo (clk, count, data_in, data_out, fifo_reset, overrun, pop, push, reset_status, wb_rst_i);

endmodule
