module uart_receiver (clk, counter_b, counter_t, enable, lcr, rda_int, rf_count, rf_data_out, rf_error_bit, rf_overrun, rf_pop, rx_lsr_mask, rx_reset, srx_pad_i, wb_rst_i);

endmodule
