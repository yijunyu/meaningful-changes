module uart_top (cts_pad_i, dcd_pad_i, dsr_pad_i, dtr_pad_o, int_o, ri_pad_i, rts_pad_o, srx_pad_i, stx_pad_o, wb_ack_o, wb_adr_i, wb_clk_i, wb_cyc_i, wb_dat_i, wb_dat_o, wb_rst_i, wb_sel_i, wb_stb_i, wb_we_i);

endmodule
