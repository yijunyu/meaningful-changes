module uart_wb (clk, re_o, wb_ack_o, wb_adr_i, wb_adr_int, wb_cyc_i, wb_dat32_o, wb_dat8_i, wb_dat8_o, wb_dat_i, wb_dat_o, wb_rst_i, wb_sel_i, wb_stb_i, wb_we_i, we_o);

endmodule
