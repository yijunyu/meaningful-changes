module uart_sync_flops (async_dat_i, clk_i, rst_i, stage1_clk_en_i, stage1_rst_i, sync_dat_o);

endmodule
