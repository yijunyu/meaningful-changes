module uart_transmitter (clk, enable, lcr, rx_lsr_mask, state, stx_pad_o, tf_count, tf_push, tx_reset, wb_dat_i, wb_rst_i);

endmodule
