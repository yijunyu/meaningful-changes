module uart_rfifo (clk, count, data_in, data_out, error_bit, fifo_reset, overrun, pop, push, reset_status, wb_rst_i);

endmodule
