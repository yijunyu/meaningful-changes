module uart_wb (clk, re_o, wb_ack_o, wb_cyc_i, wb_rst_i, wb_stb_i, wb_we_i, we_o);

endmodule
