module raminfr (a, clk, di, dpo, dpra, we);

endmodule
