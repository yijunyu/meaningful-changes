module uart_debug_if (fcr, ier, iir, lcr, lsr, mcr, msr, rf_count, rstate, tf_count, tstate, wb_adr_i, wb_dat32_o);

endmodule
