module uart_regs (clk, dtr_pad_o, enable, int_o, modem_inputs, rts_pad_o, srx_pad_i, stx_pad_o, wb_addr_i, wb_dat_i, wb_dat_o, wb_re_i, wb_rst_i, wb_we_i);

endmodule
