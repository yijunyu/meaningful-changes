module uart_transmitter (clk, enable, lcr, lsr_mask, stx_pad_o, tf_count, tf_push, tstate, tx_reset, wb_dat_i, wb_rst_i);

endmodule
